module cnn(clk,rst,data,
				data_b,
				data_w,
				result_en,
				result1,result2,result3,result4,result5,result6,result7,result8,result9,result10,result11,result12,result13,result14,result15,result16);
input clk;
input rst;
input [32-1 :0]data;
input [32*16-1 :0] data_b;
input [32*9*16 -1 :0] data_w;
output result_en;
output [32-1:0] result1,result2,result3,result4,result5,result6,result7,result8,result9,result10,result11,result12,result13,result14,result15,result16;

assign result_en = ken_1;

wire [32*9 -1 :0]data_kernel;
wire mul_en;
wire kernel_en;
reg ken_1;
get_data g1(clk,rst,data,data_kernel,mul_en,kernel_en);

always @(posedge clk)
begin
	ken_1 = kernel_en;
end

wire [31:0] mul11,mul12,mul13,mul14,mul15,mul16,mul17,mul18,mul19;
wire [31:0] mul21,mul22,mul23,mul24,mul25,mul26,mul27,mul28,mul29;
wire [31:0] mul31,mul32,mul33,mul34,mul35,mul36,mul37,mul38,mul39;
wire [31:0] mul41,mul42,mul43,mul44,mul45,mul46,mul47,mul48,mul49;
wire [31:0] mul51,mul52,mul53,mul54,mul55,mul56,mul57,mul58,mul59;
wire [31:0] mul61,mul62,mul63,mul64,mul65,mul66,mul67,mul68,mul69;
wire [31:0] mul71,mul72,mul73,mul74,mul75,mul76,mul77,mul78,mul79;
wire [31:0] mul81,mul82,mul83,mul84,mul85,mul86,mul87,mul88,mul89;
wire [31:0] mul91,mul92,mul93,mul94,mul95,mul96,mul97,mul98,mul99;
wire [31:0] mul101,mul102,mul103,mul104,mul105,mul106,mul107,mul108,mul109;
wire [31:0] mul111,mul112,mul113,mul114,mul115,mul116,mul117,mul118,mul119;
wire [31:0] mul121,mul122,mul123,mul124,mul125,mul126,mul127,mul128,mul129;
wire [31:0] mul131,mul132,mul133,mul134,mul135,mul136,mul137,mul138,mul139;
wire [31:0] mul141,mul142,mul143,mul144,mul145,mul146,mul147,mul148,mul149;
wire [31:0] mul151,mul152,mul153,mul154,mul155,mul156,mul157,mul158,mul159;
wire [31:0] mul161,mul162,mul163,mul164,mul165,mul166,mul167,mul168,mul169;

wire [31:0] add11,add12,add13,add14,add15,add16,add17,add18,add19;
wire [31:0] add21,add22,add23,add24,add25,add26,add27,add28,add29;
wire [31:0] add31,add32,add33,add34,add35,add36,add37,add38,add39;
wire [31:0] add41,add42,add43,add44,add45,add46,add47,add48,add49;
wire [31:0] add51,add52,add53,add54,add55,add56,add57,add58,add59;
wire [31:0] add61,add62,add63,add64,add65,add66,add67,add68,add69;
wire [31:0] add71,add72,add73,add74,add75,add76,add77,add78,add79;
wire [31:0] add81,add82,add83,add84,add85,add86,add87,add88,add89;
wire [31:0] add91,add92,add93,add94,add95,add96,add97,add98,add99;
wire [31:0] add101,add102,add103,add104,add105,add106,add107,add108,add109;
wire [31:0] add111,add112,add113,add114,add115,add116,add117,add118,add119;
wire [31:0] add121,add122,add123,add124,add125,add126,add127,add128,add129;
wire [31:0] add131,add132,add133,add134,add135,add136,add137,add138,add139;
wire [31:0] add141,add142,add143,add144,add145,add146,add147,add148,add149;
wire [31:0] add151,add152,add153,add154,add155,add156,add157,add158,add159;
wire [31:0] add161,add162,add163,add164,add165,add166,add167,add168,add169;

assign result1 = add19;
assign result2 = add29;
assign result3 = add39;
assign result4 = add49;
assign result5 = add59;
assign result6 = add69;
assign result7 = add79;
assign result8 = add89;
assign result9 = add99;
assign result10 = add109;
assign result11 = add119;
assign result12 = add129;
assign result13 = add139;
assign result14 = add149;
assign result15 = add159;
assign result16 = add169;

mul m11(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[31:0]),.flout_c(mul11),.round_cfg(1'b0),.en(mul_en));
mul m12(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[63:32]),.flout_c(mul12),.round_cfg(1'b0),.en(mul_en));
mul m13(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[95:64]),.flout_c(mul13),.round_cfg(1'b0),.en(mul_en));
mul m14(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[127:96]),.flout_c(mul14),.round_cfg(1'b0),.en(mul_en));
mul m15(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[159:128]),.flout_c(mul15),.round_cfg(1'b0),.en(mul_en));
mul m16(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[191:160]),.flout_c(mul16),.round_cfg(1'b0),.en(mul_en));
mul m17(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[223:192]),.flout_c(mul17),.round_cfg(1'b0),.en(mul_en));
mul m18(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[255:224]),.flout_c(mul18),.round_cfg(1'b0),.en(mul_en));
mul m19(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[287:256]),.flout_c(mul19),.round_cfg(1'b0),.en(mul_en));
mul m21(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[319:288]),.flout_c(mul21),.round_cfg(1'b0),.en(mul_en));
mul m22(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[351:320]),.flout_c(mul22),.round_cfg(1'b0),.en(mul_en));
mul m23(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[383:352]),.flout_c(mul23),.round_cfg(1'b0),.en(mul_en));
mul m24(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[415:384]),.flout_c(mul24),.round_cfg(1'b0),.en(mul_en));
mul m25(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[447:416]),.flout_c(mul25),.round_cfg(1'b0),.en(mul_en));
mul m26(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[479:448]),.flout_c(mul26),.round_cfg(1'b0),.en(mul_en));
mul m27(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[511:480]),.flout_c(mul27),.round_cfg(1'b0),.en(mul_en));
mul m28(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[543:512]),.flout_c(mul28),.round_cfg(1'b0),.en(mul_en));
mul m29(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[575:544]),.flout_c(mul29),.round_cfg(1'b0),.en(mul_en));
mul m31(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[607:576]),.flout_c(mul31),.round_cfg(1'b0),.en(mul_en));
mul m32(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[639:608]),.flout_c(mul32),.round_cfg(1'b0),.en(mul_en));
mul m33(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[671:640]),.flout_c(mul33),.round_cfg(1'b0),.en(mul_en));
mul m34(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[703:672]),.flout_c(mul34),.round_cfg(1'b0),.en(mul_en));
mul m35(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[735:704]),.flout_c(mul35),.round_cfg(1'b0),.en(mul_en));
mul m36(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[767:736]),.flout_c(mul36),.round_cfg(1'b0),.en(mul_en));
mul m37(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[799:768]),.flout_c(mul37),.round_cfg(1'b0),.en(mul_en));
mul m38(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[831:800]),.flout_c(mul38),.round_cfg(1'b0),.en(mul_en));
mul m39(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[863:832]),.flout_c(mul39),.round_cfg(1'b0),.en(mul_en));
mul m41(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[895:864]),.flout_c(mul41),.round_cfg(1'b0),.en(mul_en));
mul m42(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[927:896]),.flout_c(mul42),.round_cfg(1'b0),.en(mul_en));
mul m43(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[959:928]),.flout_c(mul43),.round_cfg(1'b0),.en(mul_en));
mul m44(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[991:960]),.flout_c(mul44),.round_cfg(1'b0),.en(mul_en));
mul m45(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[1023:992]),.flout_c(mul45),.round_cfg(1'b0),.en(mul_en));
mul m46(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[1055:1024]),.flout_c(mul46),.round_cfg(1'b0),.en(mul_en));
mul m47(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[1087:1056]),.flout_c(mul47),.round_cfg(1'b0),.en(mul_en));
mul m48(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[1119:1088]),.flout_c(mul48),.round_cfg(1'b0),.en(mul_en));
mul m49(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[1151:1120]),.flout_c(mul49),.round_cfg(1'b0),.en(mul_en));
mul m51(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[1183:1152]),.flout_c(mul51),.round_cfg(1'b0),.en(mul_en));
mul m52(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[1215:1184]),.flout_c(mul52),.round_cfg(1'b0),.en(mul_en));
mul m53(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[1247:1216]),.flout_c(mul53),.round_cfg(1'b0),.en(mul_en));
mul m54(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[1279:1248]),.flout_c(mul54),.round_cfg(1'b0),.en(mul_en));
mul m55(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[1311:1280]),.flout_c(mul55),.round_cfg(1'b0),.en(mul_en));
mul m56(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[1343:1312]),.flout_c(mul56),.round_cfg(1'b0),.en(mul_en));
mul m57(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[1375:1344]),.flout_c(mul57),.round_cfg(1'b0),.en(mul_en));
mul m58(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[1407:1376]),.flout_c(mul58),.round_cfg(1'b0),.en(mul_en));
mul m59(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[1439:1408]),.flout_c(mul59),.round_cfg(1'b0),.en(mul_en));
mul m61(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[1471:1440]),.flout_c(mul61),.round_cfg(1'b0),.en(mul_en));
mul m62(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[1503:1472]),.flout_c(mul62),.round_cfg(1'b0),.en(mul_en));
mul m63(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[1535:1504]),.flout_c(mul63),.round_cfg(1'b0),.en(mul_en));
mul m64(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[1567:1536]),.flout_c(mul64),.round_cfg(1'b0),.en(mul_en));
mul m65(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[1599:1568]),.flout_c(mul65),.round_cfg(1'b0),.en(mul_en));
mul m66(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[1631:1600]),.flout_c(mul66),.round_cfg(1'b0),.en(mul_en));
mul m67(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[1663:1632]),.flout_c(mul67),.round_cfg(1'b0),.en(mul_en));
mul m68(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[1695:1664]),.flout_c(mul68),.round_cfg(1'b0),.en(mul_en));
mul m69(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[1727:1696]),.flout_c(mul69),.round_cfg(1'b0),.en(mul_en));
mul m71(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[1759:1728]),.flout_c(mul71),.round_cfg(1'b0),.en(mul_en));
mul m72(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[1791:1760]),.flout_c(mul72),.round_cfg(1'b0),.en(mul_en));
mul m73(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[1823:1792]),.flout_c(mul73),.round_cfg(1'b0),.en(mul_en));
mul m74(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[1855:1824]),.flout_c(mul74),.round_cfg(1'b0),.en(mul_en));
mul m75(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[1887:1856]),.flout_c(mul75),.round_cfg(1'b0),.en(mul_en));
mul m76(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[1919:1888]),.flout_c(mul76),.round_cfg(1'b0),.en(mul_en));
mul m77(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[1951:1920]),.flout_c(mul77),.round_cfg(1'b0),.en(mul_en));
mul m78(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[1983:1952]),.flout_c(mul78),.round_cfg(1'b0),.en(mul_en));
mul m79(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[2015:1984]),.flout_c(mul79),.round_cfg(1'b0),.en(mul_en));
mul m81(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[2047:2016]),.flout_c(mul81),.round_cfg(1'b0),.en(mul_en));
mul m82(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[2079:2048]),.flout_c(mul82),.round_cfg(1'b0),.en(mul_en));
mul m83(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[2111:2080]),.flout_c(mul83),.round_cfg(1'b0),.en(mul_en));
mul m84(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[2143:2112]),.flout_c(mul84),.round_cfg(1'b0),.en(mul_en));
mul m85(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[2175:2144]),.flout_c(mul85),.round_cfg(1'b0),.en(mul_en));
mul m86(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[2207:2176]),.flout_c(mul86),.round_cfg(1'b0),.en(mul_en));
mul m87(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[2239:2208]),.flout_c(mul87),.round_cfg(1'b0),.en(mul_en));
mul m88(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[2271:2240]),.flout_c(mul88),.round_cfg(1'b0),.en(mul_en));
mul m89(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[2303:2272]),.flout_c(mul89),.round_cfg(1'b0),.en(mul_en));
mul m91(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[2335:2304]),.flout_c(mul91),.round_cfg(1'b0),.en(mul_en));
mul m92(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[2367:2336]),.flout_c(mul92),.round_cfg(1'b0),.en(mul_en));
mul m93(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[2399:2368]),.flout_c(mul93),.round_cfg(1'b0),.en(mul_en));
mul m94(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[2431:2400]),.flout_c(mul94),.round_cfg(1'b0),.en(mul_en));
mul m95(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[2463:2432]),.flout_c(mul95),.round_cfg(1'b0),.en(mul_en));
mul m96(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[2495:2464]),.flout_c(mul96),.round_cfg(1'b0),.en(mul_en));
mul m97(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[2527:2496]),.flout_c(mul97),.round_cfg(1'b0),.en(mul_en));
mul m98(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[2559:2528]),.flout_c(mul98),.round_cfg(1'b0),.en(mul_en));
mul m99(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[2591:2560]),.flout_c(mul99),.round_cfg(1'b0),.en(mul_en));
mul m101(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[2623:2592]),.flout_c(mul101),.round_cfg(1'b0),.en(mul_en));
mul m102(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[2655:2624]),.flout_c(mul102),.round_cfg(1'b0),.en(mul_en));
mul m103(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[2687:2656]),.flout_c(mul103),.round_cfg(1'b0),.en(mul_en));
mul m104(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[2719:2688]),.flout_c(mul104),.round_cfg(1'b0),.en(mul_en));
mul m105(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[2751:2720]),.flout_c(mul105),.round_cfg(1'b0),.en(mul_en));
mul m106(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[2783:2752]),.flout_c(mul106),.round_cfg(1'b0),.en(mul_en));
mul m107(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[2815:2784]),.flout_c(mul107),.round_cfg(1'b0),.en(mul_en));
mul m108(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[2847:2816]),.flout_c(mul108),.round_cfg(1'b0),.en(mul_en));
mul m109(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[2879:2848]),.flout_c(mul109),.round_cfg(1'b0),.en(mul_en));
mul m111(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[2911:2880]),.flout_c(mul111),.round_cfg(1'b0),.en(mul_en));
mul m112(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[2943:2912]),.flout_c(mul112),.round_cfg(1'b0),.en(mul_en));
mul m113(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[2975:2944]),.flout_c(mul113),.round_cfg(1'b0),.en(mul_en));
mul m114(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[3007:2976]),.flout_c(mul114),.round_cfg(1'b0),.en(mul_en));
mul m115(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[3039:3008]),.flout_c(mul115),.round_cfg(1'b0),.en(mul_en));
mul m116(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[3071:3040]),.flout_c(mul116),.round_cfg(1'b0),.en(mul_en));
mul m117(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[3103:3072]),.flout_c(mul117),.round_cfg(1'b0),.en(mul_en));
mul m118(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[3135:3104]),.flout_c(mul118),.round_cfg(1'b0),.en(mul_en));
mul m119(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[3167:3136]),.flout_c(mul119),.round_cfg(1'b0),.en(mul_en));
mul m121(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[3199:3168]),.flout_c(mul121),.round_cfg(1'b0),.en(mul_en));
mul m122(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[3231:3200]),.flout_c(mul122),.round_cfg(1'b0),.en(mul_en));
mul m123(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[3263:3232]),.flout_c(mul123),.round_cfg(1'b0),.en(mul_en));
mul m124(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[3295:3264]),.flout_c(mul124),.round_cfg(1'b0),.en(mul_en));
mul m125(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[3327:3296]),.flout_c(mul125),.round_cfg(1'b0),.en(mul_en));
mul m126(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[3359:3328]),.flout_c(mul126),.round_cfg(1'b0),.en(mul_en));
mul m127(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[3391:3360]),.flout_c(mul127),.round_cfg(1'b0),.en(mul_en));
mul m128(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[3423:3392]),.flout_c(mul128),.round_cfg(1'b0),.en(mul_en));
mul m129(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[3455:3424]),.flout_c(mul129),.round_cfg(1'b0),.en(mul_en));
mul m131(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[3487:3456]),.flout_c(mul131),.round_cfg(1'b0),.en(mul_en));
mul m132(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[3519:3488]),.flout_c(mul132),.round_cfg(1'b0),.en(mul_en));
mul m133(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[3551:3520]),.flout_c(mul133),.round_cfg(1'b0),.en(mul_en));
mul m134(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[3583:3552]),.flout_c(mul134),.round_cfg(1'b0),.en(mul_en));
mul m135(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[3615:3584]),.flout_c(mul135),.round_cfg(1'b0),.en(mul_en));
mul m136(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[3647:3616]),.flout_c(mul136),.round_cfg(1'b0),.en(mul_en));
mul m137(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[3679:3648]),.flout_c(mul137),.round_cfg(1'b0),.en(mul_en));
mul m138(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[3711:3680]),.flout_c(mul138),.round_cfg(1'b0),.en(mul_en));
mul m139(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[3743:3712]),.flout_c(mul139),.round_cfg(1'b0),.en(mul_en));
mul m141(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[3775:3744]),.flout_c(mul141),.round_cfg(1'b0),.en(mul_en));
mul m142(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[3807:3776]),.flout_c(mul142),.round_cfg(1'b0),.en(mul_en));
mul m143(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[3839:3808]),.flout_c(mul143),.round_cfg(1'b0),.en(mul_en));
mul m144(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[3871:3840]),.flout_c(mul144),.round_cfg(1'b0),.en(mul_en));
mul m145(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[3903:3872]),.flout_c(mul145),.round_cfg(1'b0),.en(mul_en));
mul m146(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[3935:3904]),.flout_c(mul146),.round_cfg(1'b0),.en(mul_en));
mul m147(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[3967:3936]),.flout_c(mul147),.round_cfg(1'b0),.en(mul_en));
mul m148(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[3999:3968]),.flout_c(mul148),.round_cfg(1'b0),.en(mul_en));
mul m149(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[4031:4000]),.flout_c(mul149),.round_cfg(1'b0),.en(mul_en));
mul m151(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[4063:4032]),.flout_c(mul151),.round_cfg(1'b0),.en(mul_en));
mul m152(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[4095:4064]),.flout_c(mul152),.round_cfg(1'b0),.en(mul_en));
mul m153(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[4127:4096]),.flout_c(mul153),.round_cfg(1'b0),.en(mul_en));
mul m154(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[4159:4128]),.flout_c(mul154),.round_cfg(1'b0),.en(mul_en));
mul m155(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[4191:4160]),.flout_c(mul155),.round_cfg(1'b0),.en(mul_en));
mul m156(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[4223:4192]),.flout_c(mul156),.round_cfg(1'b0),.en(mul_en));
mul m157(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[4255:4224]),.flout_c(mul157),.round_cfg(1'b0),.en(mul_en));
mul m158(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[4287:4256]),.flout_c(mul158),.round_cfg(1'b0),.en(mul_en));
mul m159(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[4319:4288]),.flout_c(mul159),.round_cfg(1'b0),.en(mul_en));
mul m161(.clk(clk),.rst(rst),.flout_a(data_kernel[31:0]),.flout_b(data_w[4351:4320]),.flout_c(mul161),.round_cfg(1'b0),.en(mul_en));
mul m162(.clk(clk),.rst(rst),.flout_a(data_kernel[63:32]),.flout_b(data_w[4383:4352]),.flout_c(mul162),.round_cfg(1'b0),.en(mul_en));
mul m163(.clk(clk),.rst(rst),.flout_a(data_kernel[95:64]),.flout_b(data_w[4415:4384]),.flout_c(mul163),.round_cfg(1'b0),.en(mul_en));
mul m164(.clk(clk),.rst(rst),.flout_a(data_kernel[127:96]),.flout_b(data_w[4447:4416]),.flout_c(mul164),.round_cfg(1'b0),.en(mul_en));
mul m165(.clk(clk),.rst(rst),.flout_a(data_kernel[159:128]),.flout_b(data_w[4479:4448]),.flout_c(mul165),.round_cfg(1'b0),.en(mul_en));
mul m166(.clk(clk),.rst(rst),.flout_a(data_kernel[191:160]),.flout_b(data_w[4511:4480]),.flout_c(mul166),.round_cfg(1'b0),.en(mul_en));
mul m167(.clk(clk),.rst(rst),.flout_a(data_kernel[223:192]),.flout_b(data_w[4543:4512]),.flout_c(mul167),.round_cfg(1'b0),.en(mul_en));
mul m168(.clk(clk),.rst(rst),.flout_a(data_kernel[255:224]),.flout_b(data_w[4575:4544]),.flout_c(mul168),.round_cfg(1'b0),.en(mul_en));
mul m169(.clk(clk),.rst(rst),.flout_a(data_kernel[287:256]),.flout_b(data_w[4607:4576]),.flout_c(mul169),.round_cfg(1'b0),.en(mul_en));


add a11(.MAIN_CLK(clk),.a(mul11),.b(mul12),.ab(add11));
add a12(.MAIN_CLK(clk),.a(add11),.b(mul13),.ab(add12));
add a13(.MAIN_CLK(clk),.a(mul14),.b(mul15),.ab(add13));
add a14(.MAIN_CLK(clk),.a(add13),.b(mul16),.ab(add14));
add a15(.MAIN_CLK(clk),.a(mul17),.b(mul18),.ab(add15));
add a16(.MAIN_CLK(clk),.a(add15),.b(mul19),.ab(add16));
add a17(.MAIN_CLK(clk),.a(add12),.b(add14),.ab(add17));
add a18(.MAIN_CLK(clk),.a(add16),.b(add17),.ab(add18));
add a19(.MAIN_CLK(clk),.a(add18),.b(data_b[31:0]),.ab(add19));
add a21(.MAIN_CLK(clk),.a(mul21),.b(mul22),.ab(add21));
add a22(.MAIN_CLK(clk),.a(add21),.b(mul23),.ab(add22));
add a23(.MAIN_CLK(clk),.a(mul24),.b(mul25),.ab(add23));
add a24(.MAIN_CLK(clk),.a(add23),.b(mul26),.ab(add24));
add a25(.MAIN_CLK(clk),.a(mul27),.b(mul28),.ab(add25));
add a26(.MAIN_CLK(clk),.a(add25),.b(mul29),.ab(add26));
add a27(.MAIN_CLK(clk),.a(add22),.b(add24),.ab(add27));
add a28(.MAIN_CLK(clk),.a(add26),.b(add27),.ab(add28));
add a29(.MAIN_CLK(clk),.a(add28),.b(data_b[63:32]),.ab(add29));
add a31(.MAIN_CLK(clk),.a(mul31),.b(mul32),.ab(add31));
add a32(.MAIN_CLK(clk),.a(add31),.b(mul33),.ab(add32));
add a33(.MAIN_CLK(clk),.a(mul34),.b(mul35),.ab(add33));
add a34(.MAIN_CLK(clk),.a(add33),.b(mul36),.ab(add34));
add a35(.MAIN_CLK(clk),.a(mul37),.b(mul38),.ab(add35));
add a36(.MAIN_CLK(clk),.a(add35),.b(mul39),.ab(add36));
add a37(.MAIN_CLK(clk),.a(add32),.b(add34),.ab(add37));
add a38(.MAIN_CLK(clk),.a(add36),.b(add37),.ab(add38));
add a39(.MAIN_CLK(clk),.a(add38),.b(data_b[95:64]),.ab(add39));
add a41(.MAIN_CLK(clk),.a(mul41),.b(mul42),.ab(add41));
add a42(.MAIN_CLK(clk),.a(add41),.b(mul43),.ab(add42));
add a43(.MAIN_CLK(clk),.a(mul44),.b(mul45),.ab(add43));
add a44(.MAIN_CLK(clk),.a(add43),.b(mul46),.ab(add44));
add a45(.MAIN_CLK(clk),.a(mul47),.b(mul48),.ab(add45));
add a46(.MAIN_CLK(clk),.a(add45),.b(mul49),.ab(add46));
add a47(.MAIN_CLK(clk),.a(add42),.b(add44),.ab(add47));
add a48(.MAIN_CLK(clk),.a(add46),.b(add47),.ab(add48));
add a49(.MAIN_CLK(clk),.a(add48),.b(data_b[127:96]),.ab(add49));
add a51(.MAIN_CLK(clk),.a(mul51),.b(mul52),.ab(add51));
add a52(.MAIN_CLK(clk),.a(add51),.b(mul53),.ab(add52));
add a53(.MAIN_CLK(clk),.a(mul54),.b(mul55),.ab(add53));
add a54(.MAIN_CLK(clk),.a(add53),.b(mul56),.ab(add54));
add a55(.MAIN_CLK(clk),.a(mul57),.b(mul58),.ab(add55));
add a56(.MAIN_CLK(clk),.a(add55),.b(mul59),.ab(add56));
add a57(.MAIN_CLK(clk),.a(add52),.b(add54),.ab(add57));
add a58(.MAIN_CLK(clk),.a(add56),.b(add57),.ab(add58));
add a59(.MAIN_CLK(clk),.a(add58),.b(data_b[159:128]),.ab(add59));
add a61(.MAIN_CLK(clk),.a(mul61),.b(mul62),.ab(add61));
add a62(.MAIN_CLK(clk),.a(add61),.b(mul63),.ab(add62));
add a63(.MAIN_CLK(clk),.a(mul64),.b(mul65),.ab(add63));
add a64(.MAIN_CLK(clk),.a(add63),.b(mul66),.ab(add64));
add a65(.MAIN_CLK(clk),.a(mul67),.b(mul68),.ab(add65));
add a66(.MAIN_CLK(clk),.a(add65),.b(mul69),.ab(add66));
add a67(.MAIN_CLK(clk),.a(add62),.b(add64),.ab(add67));
add a68(.MAIN_CLK(clk),.a(add66),.b(add67),.ab(add68));
add a69(.MAIN_CLK(clk),.a(add68),.b(data_b[191:160]),.ab(add69));
add a71(.MAIN_CLK(clk),.a(mul71),.b(mul72),.ab(add71));
add a72(.MAIN_CLK(clk),.a(add71),.b(mul73),.ab(add72));
add a73(.MAIN_CLK(clk),.a(mul74),.b(mul75),.ab(add73));
add a74(.MAIN_CLK(clk),.a(add73),.b(mul76),.ab(add74));
add a75(.MAIN_CLK(clk),.a(mul77),.b(mul78),.ab(add75));
add a76(.MAIN_CLK(clk),.a(add75),.b(mul79),.ab(add76));
add a77(.MAIN_CLK(clk),.a(add72),.b(add74),.ab(add77));
add a78(.MAIN_CLK(clk),.a(add76),.b(add77),.ab(add78));
add a79(.MAIN_CLK(clk),.a(add78),.b(data_b[223:192]),.ab(add79));
add a81(.MAIN_CLK(clk),.a(mul81),.b(mul82),.ab(add81));
add a82(.MAIN_CLK(clk),.a(add81),.b(mul83),.ab(add82));
add a83(.MAIN_CLK(clk),.a(mul84),.b(mul85),.ab(add83));
add a84(.MAIN_CLK(clk),.a(add83),.b(mul86),.ab(add84));
add a85(.MAIN_CLK(clk),.a(mul87),.b(mul88),.ab(add85));
add a86(.MAIN_CLK(clk),.a(add85),.b(mul89),.ab(add86));
add a87(.MAIN_CLK(clk),.a(add82),.b(add84),.ab(add87));
add a88(.MAIN_CLK(clk),.a(add86),.b(add87),.ab(add88));
add a89(.MAIN_CLK(clk),.a(add88),.b(data_b[255:224]),.ab(add89));
add a91(.MAIN_CLK(clk),.a(mul91),.b(mul92),.ab(add91));
add a92(.MAIN_CLK(clk),.a(add91),.b(mul93),.ab(add92));
add a93(.MAIN_CLK(clk),.a(mul94),.b(mul95),.ab(add93));
add a94(.MAIN_CLK(clk),.a(add93),.b(mul96),.ab(add94));
add a95(.MAIN_CLK(clk),.a(mul97),.b(mul98),.ab(add95));
add a96(.MAIN_CLK(clk),.a(add95),.b(mul99),.ab(add96));
add a97(.MAIN_CLK(clk),.a(add92),.b(add94),.ab(add97));
add a98(.MAIN_CLK(clk),.a(add96),.b(add97),.ab(add98));
add a99(.MAIN_CLK(clk),.a(add98),.b(data_b[287:256]),.ab(add99));
add a101(.MAIN_CLK(clk),.a(mul101),.b(mul102),.ab(add101));
add a102(.MAIN_CLK(clk),.a(add101),.b(mul103),.ab(add102));
add a103(.MAIN_CLK(clk),.a(mul104),.b(mul105),.ab(add103));
add a104(.MAIN_CLK(clk),.a(add103),.b(mul106),.ab(add104));
add a105(.MAIN_CLK(clk),.a(mul107),.b(mul108),.ab(add105));
add a106(.MAIN_CLK(clk),.a(add105),.b(mul109),.ab(add106));
add a107(.MAIN_CLK(clk),.a(add102),.b(add104),.ab(add107));
add a108(.MAIN_CLK(clk),.a(add106),.b(add107),.ab(add108));
add a109(.MAIN_CLK(clk),.a(add108),.b(data_b[319:288]),.ab(add109));
add a111(.MAIN_CLK(clk),.a(mul111),.b(mul112),.ab(add111));
add a112(.MAIN_CLK(clk),.a(add111),.b(mul113),.ab(add112));
add a113(.MAIN_CLK(clk),.a(mul114),.b(mul115),.ab(add113));
add a114(.MAIN_CLK(clk),.a(add113),.b(mul116),.ab(add114));
add a115(.MAIN_CLK(clk),.a(mul117),.b(mul118),.ab(add115));
add a116(.MAIN_CLK(clk),.a(add115),.b(mul119),.ab(add116));
add a117(.MAIN_CLK(clk),.a(add112),.b(add114),.ab(add117));
add a118(.MAIN_CLK(clk),.a(add116),.b(add117),.ab(add118));
add a119(.MAIN_CLK(clk),.a(add118),.b(data_b[351:320]),.ab(add119));
add a121(.MAIN_CLK(clk),.a(mul121),.b(mul122),.ab(add121));
add a122(.MAIN_CLK(clk),.a(add121),.b(mul123),.ab(add122));
add a123(.MAIN_CLK(clk),.a(mul124),.b(mul125),.ab(add123));
add a124(.MAIN_CLK(clk),.a(add123),.b(mul126),.ab(add124));
add a125(.MAIN_CLK(clk),.a(mul127),.b(mul128),.ab(add125));
add a126(.MAIN_CLK(clk),.a(add125),.b(mul129),.ab(add126));
add a127(.MAIN_CLK(clk),.a(add122),.b(add124),.ab(add127));
add a128(.MAIN_CLK(clk),.a(add126),.b(add127),.ab(add128));
add a129(.MAIN_CLK(clk),.a(add128),.b(data_b[383:352]),.ab(add129));
add a131(.MAIN_CLK(clk),.a(mul131),.b(mul132),.ab(add131));
add a132(.MAIN_CLK(clk),.a(add131),.b(mul133),.ab(add132));
add a133(.MAIN_CLK(clk),.a(mul134),.b(mul135),.ab(add133));
add a134(.MAIN_CLK(clk),.a(add133),.b(mul136),.ab(add134));
add a135(.MAIN_CLK(clk),.a(mul137),.b(mul138),.ab(add135));
add a136(.MAIN_CLK(clk),.a(add135),.b(mul139),.ab(add136));
add a137(.MAIN_CLK(clk),.a(add132),.b(add134),.ab(add137));
add a138(.MAIN_CLK(clk),.a(add136),.b(add137),.ab(add138));
add a139(.MAIN_CLK(clk),.a(add138),.b(data_b[415:384]),.ab(add139));
add a141(.MAIN_CLK(clk),.a(mul141),.b(mul142),.ab(add141));
add a142(.MAIN_CLK(clk),.a(add141),.b(mul143),.ab(add142));
add a143(.MAIN_CLK(clk),.a(mul144),.b(mul145),.ab(add143));
add a144(.MAIN_CLK(clk),.a(add143),.b(mul146),.ab(add144));
add a145(.MAIN_CLK(clk),.a(mul147),.b(mul148),.ab(add145));
add a146(.MAIN_CLK(clk),.a(add145),.b(mul149),.ab(add146));
add a147(.MAIN_CLK(clk),.a(add142),.b(add144),.ab(add147));
add a148(.MAIN_CLK(clk),.a(add146),.b(add147),.ab(add148));
add a149(.MAIN_CLK(clk),.a(add148),.b(data_b[447:416]),.ab(add149));
add a151(.MAIN_CLK(clk),.a(mul151),.b(mul152),.ab(add151));
add a152(.MAIN_CLK(clk),.a(add151),.b(mul153),.ab(add152));
add a153(.MAIN_CLK(clk),.a(mul154),.b(mul155),.ab(add153));
add a154(.MAIN_CLK(clk),.a(add153),.b(mul156),.ab(add154));
add a155(.MAIN_CLK(clk),.a(mul157),.b(mul158),.ab(add155));
add a156(.MAIN_CLK(clk),.a(add155),.b(mul159),.ab(add156));
add a157(.MAIN_CLK(clk),.a(add152),.b(add154),.ab(add157));
add a158(.MAIN_CLK(clk),.a(add156),.b(add157),.ab(add158));
add a159(.MAIN_CLK(clk),.a(add158),.b(data_b[479:448]),.ab(add159));
add a161(.MAIN_CLK(clk),.a(mul161),.b(mul162),.ab(add161));
add a162(.MAIN_CLK(clk),.a(add161),.b(mul163),.ab(add162));
add a163(.MAIN_CLK(clk),.a(mul164),.b(mul165),.ab(add163));
add a164(.MAIN_CLK(clk),.a(add163),.b(mul166),.ab(add164));
add a165(.MAIN_CLK(clk),.a(mul167),.b(mul168),.ab(add165));
add a166(.MAIN_CLK(clk),.a(add165),.b(mul169),.ab(add166));
add a167(.MAIN_CLK(clk),.a(add162),.b(add164),.ab(add167));
add a168(.MAIN_CLK(clk),.a(add166),.b(add167),.ab(add168));
add a169(.MAIN_CLK(clk),.a(add168),.b(data_b[511:480]),.ab(add169));

endmodule
