`timescale 1ns/1ns
module tb;

reg clk;
reg rst;
wire [31:0] data;
wire [32*16-1:0] data_b;
wire [32*9*16 -1 :0]data_w;
wire result_en;
wire [31:0] result1,result2,result3,result4,result5,result6,result7,result8,result9,result10,result11,result12,result13,result14,result15,result16;
reg [31:0] xmem [0:28*28-1];
reg [31:0] wmem [0:9*16-1];
reg [31:0] bmem [0:16-1];
reg [31:0] addr;

initial clk = 0;

always #1 clk = ~clk;
initial 
begin 
# 3000 $stop;
end
initial begin
$readmemh("E:/CASIA/SNN_RL-co/code_part/test_cnn/xhex.txt",xmem);
$readmemh("E:/CASIA/SNN_RL-co/code_part/test_cnn/wallhex.txt",wmem);
$readmemh("E:/CASIA/SNN_RL-co/code_part/test_cnn/bhex.txt",bmem);
addr = 0;
$dumpfile("tb.vcd");
$dumpvars(0,tb);
end

always @ (posedge clk)
begin 
	addr = addr + 1;
end
assign data = xmem[addr-1];
assign data_w[31:0] = wmem[0];
assign data_w[63:32] = wmem[1];
assign data_w[95:64] = wmem[2];
assign data_w[127:96] = wmem[3];
assign data_w[159:128] = wmem[4];
assign data_w[191:160] = wmem[5];
assign data_w[223:192] = wmem[6];
assign data_w[255:224] = wmem[7];
assign data_w[287:256] = wmem[8];
assign data_w[319:288] = wmem[9];
assign data_w[351:320] = wmem[10];
assign data_w[383:352] = wmem[11];
assign data_w[415:384] = wmem[12];
assign data_w[447:416] = wmem[13];
assign data_w[479:448] = wmem[14];
assign data_w[511:480] = wmem[15];
assign data_w[543:512] = wmem[16];
assign data_w[575:544] = wmem[17];
assign data_w[607:576] = wmem[18];
assign data_w[639:608] = wmem[19];
assign data_w[671:640] = wmem[20];
assign data_w[703:672] = wmem[21];
assign data_w[735:704] = wmem[22];
assign data_w[767:736] = wmem[23];
assign data_w[799:768] = wmem[24];
assign data_w[831:800] = wmem[25];
assign data_w[863:832] = wmem[26];
assign data_w[895:864] = wmem[27];
assign data_w[927:896] = wmem[28];
assign data_w[959:928] = wmem[29];
assign data_w[991:960] = wmem[30];
assign data_w[1023:992] = wmem[31];
assign data_w[1055:1024] = wmem[32];
assign data_w[1087:1056] = wmem[33];
assign data_w[1119:1088] = wmem[34];
assign data_w[1151:1120] = wmem[35];
assign data_w[1183:1152] = wmem[36];
assign data_w[1215:1184] = wmem[37];
assign data_w[1247:1216] = wmem[38];
assign data_w[1279:1248] = wmem[39];
assign data_w[1311:1280] = wmem[40];
assign data_w[1343:1312] = wmem[41];
assign data_w[1375:1344] = wmem[42];
assign data_w[1407:1376] = wmem[43];
assign data_w[1439:1408] = wmem[44];
assign data_w[1471:1440] = wmem[45];
assign data_w[1503:1472] = wmem[46];
assign data_w[1535:1504] = wmem[47];
assign data_w[1567:1536] = wmem[48];
assign data_w[1599:1568] = wmem[49];
assign data_w[1631:1600] = wmem[50];
assign data_w[1663:1632] = wmem[51];
assign data_w[1695:1664] = wmem[52];
assign data_w[1727:1696] = wmem[53];
assign data_w[1759:1728] = wmem[54];
assign data_w[1791:1760] = wmem[55];
assign data_w[1823:1792] = wmem[56];
assign data_w[1855:1824] = wmem[57];
assign data_w[1887:1856] = wmem[58];
assign data_w[1919:1888] = wmem[59];
assign data_w[1951:1920] = wmem[60];
assign data_w[1983:1952] = wmem[61];
assign data_w[2015:1984] = wmem[62];
assign data_w[2047:2016] = wmem[63];
assign data_w[2079:2048] = wmem[64];
assign data_w[2111:2080] = wmem[65];
assign data_w[2143:2112] = wmem[66];
assign data_w[2175:2144] = wmem[67];
assign data_w[2207:2176] = wmem[68];
assign data_w[2239:2208] = wmem[69];
assign data_w[2271:2240] = wmem[70];
assign data_w[2303:2272] = wmem[71];
assign data_w[2335:2304] = wmem[72];
assign data_w[2367:2336] = wmem[73];
assign data_w[2399:2368] = wmem[74];
assign data_w[2431:2400] = wmem[75];
assign data_w[2463:2432] = wmem[76];
assign data_w[2495:2464] = wmem[77];
assign data_w[2527:2496] = wmem[78];
assign data_w[2559:2528] = wmem[79];
assign data_w[2591:2560] = wmem[80];
assign data_w[2623:2592] = wmem[81];
assign data_w[2655:2624] = wmem[82];
assign data_w[2687:2656] = wmem[83];
assign data_w[2719:2688] = wmem[84];
assign data_w[2751:2720] = wmem[85];
assign data_w[2783:2752] = wmem[86];
assign data_w[2815:2784] = wmem[87];
assign data_w[2847:2816] = wmem[88];
assign data_w[2879:2848] = wmem[89];
assign data_w[2911:2880] = wmem[90];
assign data_w[2943:2912] = wmem[91];
assign data_w[2975:2944] = wmem[92];
assign data_w[3007:2976] = wmem[93];
assign data_w[3039:3008] = wmem[94];
assign data_w[3071:3040] = wmem[95];
assign data_w[3103:3072] = wmem[96];
assign data_w[3135:3104] = wmem[97];
assign data_w[3167:3136] = wmem[98];
assign data_w[3199:3168] = wmem[99];
assign data_w[3231:3200] = wmem[100];
assign data_w[3263:3232] = wmem[101];
assign data_w[3295:3264] = wmem[102];
assign data_w[3327:3296] = wmem[103];
assign data_w[3359:3328] = wmem[104];
assign data_w[3391:3360] = wmem[105];
assign data_w[3423:3392] = wmem[106];
assign data_w[3455:3424] = wmem[107];
assign data_w[3487:3456] = wmem[108];
assign data_w[3519:3488] = wmem[109];
assign data_w[3551:3520] = wmem[110];
assign data_w[3583:3552] = wmem[111];
assign data_w[3615:3584] = wmem[112];
assign data_w[3647:3616] = wmem[113];
assign data_w[3679:3648] = wmem[114];
assign data_w[3711:3680] = wmem[115];
assign data_w[3743:3712] = wmem[116];
assign data_w[3775:3744] = wmem[117];
assign data_w[3807:3776] = wmem[118];
assign data_w[3839:3808] = wmem[119];
assign data_w[3871:3840] = wmem[120];
assign data_w[3903:3872] = wmem[121];
assign data_w[3935:3904] = wmem[122];
assign data_w[3967:3936] = wmem[123];
assign data_w[3999:3968] = wmem[124];
assign data_w[4031:4000] = wmem[125];
assign data_w[4063:4032] = wmem[126];
assign data_w[4095:4064] = wmem[127];
assign data_w[4127:4096] = wmem[128];
assign data_w[4159:4128] = wmem[129];
assign data_w[4191:4160] = wmem[130];
assign data_w[4223:4192] = wmem[131];
assign data_w[4255:4224] = wmem[132];
assign data_w[4287:4256] = wmem[133];
assign data_w[4319:4288] = wmem[134];
assign data_w[4351:4320] = wmem[135];
assign data_w[4383:4352] = wmem[136];
assign data_w[4415:4384] = wmem[137];
assign data_w[4447:4416] = wmem[138];
assign data_w[4479:4448] = wmem[139];
assign data_w[4511:4480] = wmem[140];
assign data_w[4543:4512] = wmem[141];
assign data_w[4575:4544] = wmem[142];
assign data_w[4607:4576] = wmem[143];

assign data_b[31:0] = bmem[0];
assign data_b[63:32] = bmem[1];
assign data_b[95:64] = bmem[2];
assign data_b[127:96] = bmem[3];
assign data_b[159:128] = bmem[4];
assign data_b[191:160] = bmem[5];
assign data_b[223:192] = bmem[6];
assign data_b[255:224] = bmem[7];
assign data_b[287:256] = bmem[8];
assign data_b[319:288] = bmem[9];
assign data_b[351:320] = bmem[10];
assign data_b[383:352] = bmem[11];
assign data_b[415:384] = bmem[12];
assign data_b[447:416] = bmem[13];
assign data_b[479:448] = bmem[14];
assign data_b[511:480] = bmem[15];


cnn c1(clk,rst,data,data_b,data_w,result_en,result1,result2,result3,result4,result5,result6,result7,result8,result9,result10,result11,result12,result13,result14,result15,result16);

endmodule 